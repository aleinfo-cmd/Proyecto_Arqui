`timescale 1ns/1ns
module AND (
    input A,
    input B,
    output salida
);
    
assign salida = A && B;

endmodule